// ELEX 7660 Project - HDMI
// Main module to test the usage of the HDMI module
// Michael Andrews 2021/03/29

`define DIVISOR 10
`define TESTNUM 10

module AV_Top ( output [2:0] TMDSp, TMDSn, 
				output TMDSp_clock, TMDSn_clock, clk_68, rgb_clk,
				input reset_n, FPGA_CLK1_50, 

                //ADC signals, must be pin planned in top level module
                (* altera_attribute = "-name WEAK_PULL_UP_RESISTOR ON" *)
	            output ADC_CONVST, ADC_SCK, ADC_SDI,
	            input ADC_SDO
);
					
	logic clk, valid; // clock
    logic [1:0] redMag, blueMag, greenMag, whiteMag;
    logic [7:0] clkCount;
    //dft output
    logic signed [31:0] mag0;
    logic signed [31:0] mag1;
    logic signed [31:0] mag2;
    logic signed [31:0] mag3;
    logic [2:0] adc_channel = 'd0; //ADC channel to sample

    pll pll0 ( .inclk0(FPGA_CLK1_50), .c0(clk) ) ;
	HDMI HDMI_0 ( .pixelClk(clk), .redMag, .blueMag, .greenMag, .whiteMag, .TMDSp, .TMDSn, .TMDSp_clock, .TMDSn_clock ) ;
    dft dft_0 ( .clk(clk_68), .reset_n, .valid, .mag0, .mag1, .mag2, .mag3 , .ADC_CONVST, .ADC_SCK, .ADC_SDI, .ADC_SDO, .adc_channel ) ;

    always_ff @( posedge valid ) begin
        whiteMag <= mag0[13:12];
        blueMag <= mag1[11:10];
        greenMag <= mag2[12:11];
        redMag <= mag3[11:10];
    end
    

    /*always_comb begin
        //Testing block
        if (magX[0] < `TESTNUM) begin
            rgb_clk = 0;
        end
        else begin
            rgb_clk = 1;
        end
    end*/

    //Clock divider to create a 68kHz clock for the ADC
    always_ff @(posedge clk) begin
        if (clkCount == 'd183) begin
            clkCount <= 'd0;
            clk_68 <= ~clk_68;
        end
        else
            clkCount <= clkCount + 1;
    end
endmodule

// megafunction wizard: %ALTPLL%
// ...
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
// ...

module pll ( inclk0, c0);

        input     inclk0;
        output    c0;

        wire [0:0] sub_wire2 = 1'h0;
        wire [4:0] sub_wire3;
        wire  sub_wire0 = inclk0;
        wire [1:0] sub_wire1 = {sub_wire2, sub_wire0};
        wire [0:0] sub_wire4 = sub_wire3[0:0];
        wire  c0 = sub_wire4;

        altpll altpll_component ( .inclk (sub_wire1), .clk
          (sub_wire3), .activeclock (), .areset (1'b0), .clkbad
          (), .clkena ({6{1'b1}}), .clkloss (), .clkswitch
          (1'b0), .configupdate (1'b0), .enable0 (), .enable1 (),
          .extclk (), .extclkena ({4{1'b1}}), .fbin (1'b1),
          .fbmimicbidir (), .fbout (), .fref (), .icdrclk (),
          .locked (), .pfdena (1'b1), .phasecounterselect
          ({4{1'b1}}), .phasedone (), .phasestep (1'b1),
          .phaseupdown (1'b1), .pllena (1'b1), .scanaclr (1'b0),
          .scanclk (1'b0), .scanclkena (1'b1), .scandata (1'b0),
          .scandataout (), .scandone (), .scanread (1'b0),
          .scanwrite (1'b0), .sclkout0 (), .sclkout1 (),
          .vcooverrange (), .vcounderrange ());

        defparam
                altpll_component.bandwidth_type = "AUTO",
                altpll_component.clk0_divide_by = 2,
                altpll_component.clk0_duty_cycle = 50,
                altpll_component.clk0_multiply_by = 1,
                altpll_component.clk0_phase_shift = "0",
                altpll_component.compensate_clock = "CLK0",
                altpll_component.inclk0_input_frequency = 20000,
                altpll_component.intended_device_family = "Cyclone IV E",
                altpll_component.lpm_hint = "CBX_MODULE_PREFIX=lab1clk",
                altpll_component.lpm_type = "altpll",
                altpll_component.operation_mode = "NORMAL",
                altpll_component.pll_type = "AUTO",
                altpll_component.port_activeclock = "PORT_UNUSED",
                altpll_component.port_areset = "PORT_UNUSED",
                altpll_component.port_clkbad0 = "PORT_UNUSED",
                altpll_component.port_clkbad1 = "PORT_UNUSED",
                altpll_component.port_clkloss = "PORT_UNUSED",
                altpll_component.port_clkswitch = "PORT_UNUSED",
                altpll_component.port_configupdate = "PORT_UNUSED",
                altpll_component.port_fbin = "PORT_UNUSED",
                altpll_component.port_inclk0 = "PORT_USED",
                altpll_component.port_inclk1 = "PORT_UNUSED",
                altpll_component.port_locked = "PORT_UNUSED",
                altpll_component.port_pfdena = "PORT_UNUSED",
                altpll_component.port_phasecounterselect = "PORT_UNUSED",
                altpll_component.port_phasedone = "PORT_UNUSED",
                altpll_component.port_phasestep = "PORT_UNUSED",
                altpll_component.port_phaseupdown = "PORT_UNUSED",
                altpll_component.port_pllena = "PORT_UNUSED",
                altpll_component.port_scanaclr = "PORT_UNUSED",
                altpll_component.port_scanclk = "PORT_UNUSED",
                altpll_component.port_scanclkena = "PORT_UNUSED",
                altpll_component.port_scandata = "PORT_UNUSED",
                altpll_component.port_scandataout = "PORT_UNUSED",
                altpll_component.port_scandone = "PORT_UNUSED",
                altpll_component.port_scanread = "PORT_UNUSED",
                altpll_component.port_scanwrite = "PORT_UNUSED",
                altpll_component.port_clk0 = "PORT_USED",
                altpll_component.port_clk1 = "PORT_UNUSED",
                altpll_component.port_clk2 = "PORT_UNUSED",
                altpll_component.port_clk3 = "PORT_UNUSED",
                altpll_component.port_clk4 = "PORT_UNUSED",
                altpll_component.port_clk5 = "PORT_UNUSED",
                altpll_component.port_clkena0 = "PORT_UNUSED",
                altpll_component.port_clkena1 = "PORT_UNUSED",
                altpll_component.port_clkena2 = "PORT_UNUSED",
                altpll_component.port_clkena3 = "PORT_UNUSED",
                altpll_component.port_clkena4 = "PORT_UNUSED",
                altpll_component.port_clkena5 = "PORT_UNUSED",
                altpll_component.port_extclk0 = "PORT_UNUSED",
                altpll_component.port_extclk1 = "PORT_UNUSED",
                altpll_component.port_extclk2 = "PORT_UNUSED",
                altpll_component.port_extclk3 = "PORT_UNUSED",
                altpll_component.width_clock = 5;


endmodule